library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.pkg_axi.all;

entity zynq_ps_wrap is
    port (
        DDR_addr          : inout std_logic_vector(14 downto 0);
        DDR_ba            : inout std_logic_vector(2 downto 0);
        DDR_cas_n         : inout std_logic;
        DDR_ck_n          : inout std_logic;
        DDR_ck_p          : inout std_logic;
        DDR_cke           : inout std_logic;
        DDR_cs_n          : inout std_logic;
        DDR_dm            : inout std_logic_vector(3 downto 0);
        DDR_dq            : inout std_logic_vector(31 downto 0);
        DDR_dqs_n         : inout std_logic_vector(3 downto 0);
        DDR_dqs_p         : inout std_logic_vector(3 downto 0);
        DDR_odt           : inout std_logic;
        DDR_ras_n         : inout std_logic;
        DDR_reset_n       : inout std_logic;
        DDR_we_n          : inout std_logic;
        FIXED_IO_ddr_vrn  : inout std_logic;
        FIXED_IO_ddr_vrp  : inout std_logic;
        FIXED_IO_mio      : inout std_logic_vector(53 downto 0);
        FIXED_IO_ps_clk   : inout std_logic;
        FIXED_IO_ps_porb  : inout std_logic;
        FIXED_IO_ps_srstb : inout std_logic;
        REF_CLK           : out   std_logic;
        REF_RST           : out   std_logic;
        ACLK              : out   std_logic;
        ARESET            : out   std_logic;
        M_AXI_REG0_OUT    : out   axi4lite_mout_sin;
        M_AXI_REG0_IN     : in    axi4lite_min_sout;
        M_AXI_REG1_OUT    : out   axi4lite_mout_sin;
        M_AXI_REG1_IN     : in    axi4lite_min_sout;
        S_AXI_DRAM0_OUT   : out   axi4_min_sout;
        S_AXI_DRAM0_IN    : in    axi4_mout_sin;
        S_AXI_DRAM1_OUT   : out   axi4_min_sout;
        S_AXI_DRAM1_IN    : in    axi4_mout_sin;
        S_AXI_DRAM2_OUT   : out   axi4_min_sout;
        S_AXI_DRAM2_IN    : in    axi4_mout_sin;
        S_AXI_DRAM3_OUT   : out   axi4_min_sout;
        S_AXI_DRAM3_IN    : in    axi4_mout_sin
        );
end zynq_ps_wrap;

architecture structural of zynq_ps_wrap is

    signal REF_CLK_int : std_logic;
    signal REF_ARST    : std_logic;

begin

    rst_ref_sync : entity work.rst_synchro
        generic map (
            rst_in_active_high  => true,  -- boolean               := true;
            rst_out_active_high => true,  -- boolean               := true;
            rst_out_min_cycles  => 8      -- integer range 3 to 10 := 4
            )
        port map (
            arst => REF_ARST,             -- in  std_logic;        -- captured asynchronously
            clk  => REF_CLK_int,          -- in  std_logic;
            rst  => REF_RST               -- out std_logic         -- fully synchronous
            );

    REF_CLK <= REF_CLK_int;

    zynq_ps_wrapper_inst : entity work.zynq_ps_wrapper
        port map (
            DDR_addr             => DDR_addr,                 -- inout std_logic_vector(14 downto 0);
            DDR_ba               => DDR_ba,                   -- inout std_logic_vector(2 downto 0);
            DDR_cas_n            => DDR_cas_n,                -- inout std_logic;
            DDR_ck_n             => DDR_ck_n,                 -- inout std_logic;
            DDR_ck_p             => DDR_ck_p,                 -- inout std_logic;
            DDR_cke              => DDR_cke,                  -- inout std_logic;
            DDR_cs_n             => DDR_cs_n,                 -- inout std_logic;
            DDR_dm               => DDR_dm,                   -- inout std_logic_vector(3 downto 0);
            DDR_dq               => DDR_dq,                   -- inout std_logic_vector(31 downto 0);
            DDR_dqs_n            => DDR_dqs_n,                -- inout std_logic_vector(3 downto 0);
            DDR_dqs_p            => DDR_dqs_p,                -- inout std_logic_vector(3 downto 0);
            DDR_odt              => DDR_odt,                  -- inout std_logic;
            DDR_ras_n            => DDR_ras_n,                -- inout std_logic;
            DDR_reset_n          => DDR_reset_n,              -- inout std_logic;
            DDR_we_n             => DDR_we_n,                 -- inout std_logic;
            FIXED_IO_ddr_vrn     => FIXED_IO_ddr_vrn,         -- inout std_logic;
            FIXED_IO_ddr_vrp     => FIXED_IO_ddr_vrp,         -- inout std_logic;
            FIXED_IO_mio         => FIXED_IO_mio,             -- inout std_logic_vector(53 downto 0);
            FIXED_IO_ps_clk      => FIXED_IO_ps_clk,          -- inout std_logic;
            FIXED_IO_ps_porb     => FIXED_IO_ps_porb,         -- inout std_logic;
            FIXED_IO_ps_srstb    => FIXED_IO_ps_srstb,        -- inout std_logic;
            REF_CLK              => REF_CLK_int,              -- out   std_logic;
            REF_RST(0)           => REF_ARST,                 -- out   std_logic;
            ACLK                 => ACLK,                     -- out   std_logic;
            ARESET(0)            => ARESET,                   -- out   std_logic_vector(0 to 0);
            M_AXI_REG0_arready   => M_AXI_REG0_IN.arready,    -- in    std_logic;
            M_AXI_REG0_awready   => M_AXI_REG0_IN.awready,    -- in    std_logic;
            M_AXI_REG0_bresp     => M_AXI_REG0_IN.bresp,      -- in    std_logic_vector(1 downto 0);
            M_AXI_REG0_bvalid    => M_AXI_REG0_IN.bvalid,     -- in    std_logic;
            M_AXI_REG0_rdata     => M_AXI_REG0_IN.rdata,      -- in    std_logic_vector(31 downto 0);
            M_AXI_REG0_rresp     => M_AXI_REG0_IN.rresp,      -- in    std_logic_vector(1 downto 0);
            M_AXI_REG0_rvalid    => M_AXI_REG0_IN.rvalid,     -- in    std_logic;
            M_AXI_REG0_wready    => M_AXI_REG0_IN.wready,     -- in    std_logic;
            M_AXI_REG0_araddr    => M_AXI_REG0_OUT.araddr,    -- out   std_logic_vector(31 downto 0);
            M_AXI_REG0_arprot    => M_AXI_REG0_OUT.arprot,    -- out   std_logic_vector(2 downto 0);
            M_AXI_REG0_arvalid   => M_AXI_REG0_OUT.arvalid,   -- out   std_logic;
            M_AXI_REG0_awaddr    => M_AXI_REG0_OUT.awaddr,    -- out   std_logic_vector(31 downto 0);
            M_AXI_REG0_awprot    => M_AXI_REG0_OUT.awprot,    -- out   std_logic_vector(2 downto 0);
            M_AXI_REG0_awvalid   => M_AXI_REG0_OUT.awvalid,   -- out   std_logic;
            M_AXI_REG0_bready    => M_AXI_REG0_OUT.bready,    -- out   std_logic;
            M_AXI_REG0_rready    => M_AXI_REG0_OUT.rready,    -- out   std_logic;
            M_AXI_REG0_wdata     => M_AXI_REG0_OUT.wdata,     -- out   std_logic_vector(31 downto 0);
            M_AXI_REG0_wstrb     => M_AXI_REG0_OUT.wstrb,     -- out   std_logic_vector(3 downto 0);
            M_AXI_REG0_wvalid    => M_AXI_REG0_OUT.wvalid,    -- out   std_logic;
            M_AXI_REG1_arready   => M_AXI_REG1_IN.arready,    -- in    std_logic;
            M_AXI_REG1_awready   => M_AXI_REG1_IN.awready,    -- in    std_logic;
            M_AXI_REG1_bresp     => M_AXI_REG1_IN.bresp,      -- in    std_logic_vector(1 downto 0);
            M_AXI_REG1_bvalid    => M_AXI_REG1_IN.bvalid,     -- in    std_logic;
            M_AXI_REG1_rdata     => M_AXI_REG1_IN.rdata,      -- in    std_logic_vector(31 downto 0);
            M_AXI_REG1_rresp     => M_AXI_REG1_IN.rresp,      -- in    std_logic_vector(1 downto 0);
            M_AXI_REG1_rvalid    => M_AXI_REG1_IN.rvalid,     -- in    std_logic;
            M_AXI_REG1_wready    => M_AXI_REG1_IN.wready,     -- in    std_logic;
            M_AXI_REG1_araddr    => M_AXI_REG1_OUT.araddr,    -- out   std_logic_vector(31 downto 0);
            M_AXI_REG1_arprot    => M_AXI_REG1_OUT.arprot,    -- out   std_logic_vector(2 downto 0);
            M_AXI_REG1_arvalid   => M_AXI_REG1_OUT.arvalid,   -- out   std_logic;
            M_AXI_REG1_awaddr    => M_AXI_REG1_OUT.awaddr,    -- out   std_logic_vector(31 downto 0);
            M_AXI_REG1_awprot    => M_AXI_REG1_OUT.awprot,    -- out   std_logic_vector(2 downto 0);
            M_AXI_REG1_awvalid   => M_AXI_REG1_OUT.awvalid,   -- out   std_logic;
            M_AXI_REG1_bready    => M_AXI_REG1_OUT.bready,    -- out   std_logic;
            M_AXI_REG1_rready    => M_AXI_REG1_OUT.rready,    -- out   std_logic;
            M_AXI_REG1_wdata     => M_AXI_REG1_OUT.wdata,     -- out   std_logic_vector(31 downto 0);
            M_AXI_REG1_wstrb     => M_AXI_REG1_OUT.wstrb,     -- out   std_logic_vector(3 downto 0);
            M_AXI_REG1_wvalid    => M_AXI_REG1_OUT.wvalid,    -- out   std_logic;
            S_AXI_DRAM0_araddr   => S_AXI_DRAM0_IN.araddr,    -- in    std_logic_vector(31 downto 0);
            S_AXI_DRAM0_arburst  => S_AXI_DRAM0_IN.arburst,   -- in    std_logic_vector(1 downto 0);
            S_AXI_DRAM0_arcache  => S_AXI_DRAM0_IN.arcache,   -- in    std_logic_vector(3 downto 0);
            S_AXI_DRAM0_arlen    => S_AXI_DRAM0_IN.arlen,     -- in    std_logic_vector(7 downto 0);
            S_AXI_DRAM0_arlock   => S_AXI_DRAM0_IN.arlock,    -- in    std_logic_vector(0 to 0);
            S_AXI_DRAM0_arprot   => S_AXI_DRAM0_IN.arprot,    -- in    std_logic_vector(2 downto 0);
            S_AXI_DRAM0_arqos    => S_AXI_DRAM0_IN.arqos,     -- in    std_logic_vector(3 downto 0);
            S_AXI_DRAM0_arregion => S_AXI_DRAM0_IN.arregion,  -- in    std_logic_vector(3 downto 0);
            S_AXI_DRAM0_arsize   => S_AXI_DRAM0_IN.arsize,    -- in    std_logic_vector(2 downto 0);
            S_AXI_DRAM0_arvalid  => S_AXI_DRAM0_IN.arvalid,   -- in    std_logic;
            S_AXI_DRAM0_awaddr   => S_AXI_DRAM0_IN.awaddr,    -- in    std_logic_vector(31 downto 0);
            S_AXI_DRAM0_awburst  => S_AXI_DRAM0_IN.awburst,   -- in    std_logic_vector(1 downto 0);
            S_AXI_DRAM0_awcache  => S_AXI_DRAM0_IN.awcache,   -- in    std_logic_vector(3 downto 0);
            S_AXI_DRAM0_awlen    => S_AXI_DRAM0_IN.awlen,     -- in    std_logic_vector(7 downto 0);
            S_AXI_DRAM0_awlock   => S_AXI_DRAM0_IN.awlock,    -- in    std_logic_vector(0 to 0);
            S_AXI_DRAM0_awprot   => S_AXI_DRAM0_IN.awprot,    -- in    std_logic_vector(2 downto 0);
            S_AXI_DRAM0_awqos    => S_AXI_DRAM0_IN.awqos,     -- in    std_logic_vector(3 downto 0);
            S_AXI_DRAM0_awregion => S_AXI_DRAM0_IN.awregion,  -- in    std_logic_vector(3 downto 0);
            S_AXI_DRAM0_awsize   => S_AXI_DRAM0_IN.awsize,    -- in    std_logic_vector(2 downto 0);
            S_AXI_DRAM0_awvalid  => S_AXI_DRAM0_IN.awvalid,   -- in    std_logic;
            S_AXI_DRAM0_bready   => S_AXI_DRAM0_IN.bready,    -- in    std_logic;
            S_AXI_DRAM0_rready   => S_AXI_DRAM0_IN.rready,    -- in    std_logic;
            S_AXI_DRAM0_wdata    => S_AXI_DRAM0_IN.wdata,     -- in    std_logic_vector(63 downto 0);
            S_AXI_DRAM0_wlast    => S_AXI_DRAM0_IN.wlast,     -- in    std_logic;
            S_AXI_DRAM0_wstrb    => S_AXI_DRAM0_IN.wstrb,     -- in    std_logic_vector(7 downto 0);
            S_AXI_DRAM0_wvalid   => S_AXI_DRAM0_IN.wvalid,    -- in    std_logic;
            S_AXI_DRAM0_arready  => S_AXI_DRAM0_OUT.arready,  -- out   std_logic;
            S_AXI_DRAM0_awready  => S_AXI_DRAM0_OUT.awready,  -- out   std_logic;
            S_AXI_DRAM0_bresp    => S_AXI_DRAM0_OUT.bresp,    -- out   std_logic_vector(1 downto 0);
            S_AXI_DRAM0_bvalid   => S_AXI_DRAM0_OUT.bvalid,   -- out   std_logic;
            S_AXI_DRAM0_rdata    => S_AXI_DRAM0_OUT.rdata,    -- out   std_logic_vector(63 downto 0);
            S_AXI_DRAM0_rlast    => S_AXI_DRAM0_OUT.rlast,    -- out   std_logic;
            S_AXI_DRAM0_rresp    => S_AXI_DRAM0_OUT.rresp,    -- out   std_logic_vector(1 downto 0);
            S_AXI_DRAM0_rvalid   => S_AXI_DRAM0_OUT.rvalid,   -- out   std_logic;
            S_AXI_DRAM0_wready   => S_AXI_DRAM0_OUT.wready,   -- out   std_logic;
            S_AXI_DRAM1_araddr   => S_AXI_DRAM1_IN.araddr,    -- in    std_logic_vector(31 downto 0);
            S_AXI_DRAM1_arburst  => S_AXI_DRAM1_IN.arburst,   -- in    std_logic_vector(1 downto 0);
            S_AXI_DRAM1_arcache  => S_AXI_DRAM1_IN.arcache,   -- in    std_logic_vector(3 downto 0);
            S_AXI_DRAM1_arlen    => S_AXI_DRAM1_IN.arlen,     -- in    std_logic_vector(7 downto 0);
            S_AXI_DRAM1_arlock   => S_AXI_DRAM1_IN.arlock,    -- in    std_logic_vector(0 to 0);
            S_AXI_DRAM1_arprot   => S_AXI_DRAM1_IN.arprot,    -- in    std_logic_vector(2 downto 0);
            S_AXI_DRAM1_arqos    => S_AXI_DRAM1_IN.arqos,     -- in    std_logic_vector(3 downto 0);
            S_AXI_DRAM1_arregion => S_AXI_DRAM1_IN.arregion,  -- in    std_logic_vector(3 downto 0);
            S_AXI_DRAM1_arsize   => S_AXI_DRAM1_IN.arsize,    -- in    std_logic_vector(2 downto 0);
            S_AXI_DRAM1_arvalid  => S_AXI_DRAM1_IN.arvalid,   -- in    std_logic;
            S_AXI_DRAM1_awaddr   => S_AXI_DRAM1_IN.awaddr,    -- in    std_logic_vector(31 downto 0);
            S_AXI_DRAM1_awburst  => S_AXI_DRAM1_IN.awburst,   -- in    std_logic_vector(1 downto 0);
            S_AXI_DRAM1_awcache  => S_AXI_DRAM1_IN.awcache,   -- in    std_logic_vector(3 downto 0);
            S_AXI_DRAM1_awlen    => S_AXI_DRAM1_IN.awlen,     -- in    std_logic_vector(7 downto 0);
            S_AXI_DRAM1_awlock   => S_AXI_DRAM1_IN.awlock,    -- in    std_logic_vector(0 to 0);
            S_AXI_DRAM1_awprot   => S_AXI_DRAM1_IN.awprot,    -- in    std_logic_vector(2 downto 0);
            S_AXI_DRAM1_awqos    => S_AXI_DRAM1_IN.awqos,     -- in    std_logic_vector(3 downto 0);
            S_AXI_DRAM1_awregion => S_AXI_DRAM1_IN.awregion,  -- in    std_logic_vector(3 downto 0);
            S_AXI_DRAM1_awsize   => S_AXI_DRAM1_IN.awsize,    -- in    std_logic_vector(2 downto 0);
            S_AXI_DRAM1_awvalid  => S_AXI_DRAM1_IN.awvalid,   -- in    std_logic;
            S_AXI_DRAM1_bready   => S_AXI_DRAM1_IN.bready,    -- in    std_logic;
            S_AXI_DRAM1_rready   => S_AXI_DRAM1_IN.rready,    -- in    std_logic;
            S_AXI_DRAM1_wdata    => S_AXI_DRAM1_IN.wdata,     -- in    std_logic_vector(63 downto 0);
            S_AXI_DRAM1_wlast    => S_AXI_DRAM1_IN.wlast,     -- in    std_logic;
            S_AXI_DRAM1_wstrb    => S_AXI_DRAM1_IN.wstrb,     -- in    std_logic_vector(7 downto 0);
            S_AXI_DRAM1_wvalid   => S_AXI_DRAM1_IN.wvalid,    -- in    std_logic;
            S_AXI_DRAM1_arready  => S_AXI_DRAM1_OUT.arready,  -- out   std_logic;
            S_AXI_DRAM1_awready  => S_AXI_DRAM1_OUT.awready,  -- out   std_logic;
            S_AXI_DRAM1_bresp    => S_AXI_DRAM1_OUT.bresp,    -- out   std_logic_vector(1 downto 0);
            S_AXI_DRAM1_bvalid   => S_AXI_DRAM1_OUT.bvalid,   -- out   std_logic;
            S_AXI_DRAM1_rdata    => S_AXI_DRAM1_OUT.rdata,    -- out   std_logic_vector(63 downto 0);
            S_AXI_DRAM1_rlast    => S_AXI_DRAM1_OUT.rlast,    -- out   std_logic;
            S_AXI_DRAM1_rresp    => S_AXI_DRAM1_OUT.rresp,    -- out   std_logic_vector(1 downto 0);
            S_AXI_DRAM1_rvalid   => S_AXI_DRAM1_OUT.rvalid,   -- out   std_logic;
            S_AXI_DRAM1_wready   => S_AXI_DRAM1_OUT.wready,   -- out   std_logic;
            S_AXI_DRAM2_araddr   => S_AXI_DRAM2_IN.araddr,    -- in    std_logic_vector(31 downto 0);
            S_AXI_DRAM2_arburst  => S_AXI_DRAM2_IN.arburst,   -- in    std_logic_vector(1 downto 0);
            S_AXI_DRAM2_arcache  => S_AXI_DRAM2_IN.arcache,   -- in    std_logic_vector(3 downto 0);
            S_AXI_DRAM2_arlen    => S_AXI_DRAM2_IN.arlen,     -- in    std_logic_vector(7 downto 0);
            S_AXI_DRAM2_arlock   => S_AXI_DRAM2_IN.arlock,    -- in    std_logic_vector(0 to 0);
            S_AXI_DRAM2_arprot   => S_AXI_DRAM2_IN.arprot,    -- in    std_logic_vector(2 downto 0);
            S_AXI_DRAM2_arqos    => S_AXI_DRAM2_IN.arqos,     -- in    std_logic_vector(3 downto 0);
            S_AXI_DRAM2_arregion => S_AXI_DRAM2_IN.arregion,  -- in    std_logic_vector(3 downto 0);
            S_AXI_DRAM2_arsize   => S_AXI_DRAM2_IN.arsize,    -- in    std_logic_vector(2 downto 0);
            S_AXI_DRAM2_arvalid  => S_AXI_DRAM2_IN.arvalid,   -- in    std_logic;
            S_AXI_DRAM2_awaddr   => S_AXI_DRAM2_IN.awaddr,    -- in    std_logic_vector(31 downto 0);
            S_AXI_DRAM2_awburst  => S_AXI_DRAM2_IN.awburst,   -- in    std_logic_vector(1 downto 0);
            S_AXI_DRAM2_awcache  => S_AXI_DRAM2_IN.awcache,   -- in    std_logic_vector(3 downto 0);
            S_AXI_DRAM2_awlen    => S_AXI_DRAM2_IN.awlen,     -- in    std_logic_vector(7 downto 0);
            S_AXI_DRAM2_awlock   => S_AXI_DRAM2_IN.awlock,    -- in    std_logic_vector(0 to 0);
            S_AXI_DRAM2_awprot   => S_AXI_DRAM2_IN.awprot,    -- in    std_logic_vector(2 downto 0);
            S_AXI_DRAM2_awqos    => S_AXI_DRAM2_IN.awqos,     -- in    std_logic_vector(3 downto 0);
            S_AXI_DRAM2_awregion => S_AXI_DRAM2_IN.awregion,  -- in    std_logic_vector(3 downto 0);
            S_AXI_DRAM2_awsize   => S_AXI_DRAM2_IN.awsize,    -- in    std_logic_vector(2 downto 0);
            S_AXI_DRAM2_awvalid  => S_AXI_DRAM2_IN.awvalid,   -- in    std_logic;
            S_AXI_DRAM2_bready   => S_AXI_DRAM2_IN.bready,    -- in    std_logic;
            S_AXI_DRAM2_rready   => S_AXI_DRAM2_IN.rready,    -- in    std_logic;
            S_AXI_DRAM2_wdata    => S_AXI_DRAM2_IN.wdata,     -- in    std_logic_vector(63 downto 0);
            S_AXI_DRAM2_wlast    => S_AXI_DRAM2_IN.wlast,     -- in    std_logic;
            S_AXI_DRAM2_wstrb    => S_AXI_DRAM2_IN.wstrb,     -- in    std_logic_vector(7 downto 0);
            S_AXI_DRAM2_wvalid   => S_AXI_DRAM2_IN.wvalid,    -- in    std_logic;
            S_AXI_DRAM2_arready  => S_AXI_DRAM2_OUT.arready,  -- out   std_logic;
            S_AXI_DRAM2_awready  => S_AXI_DRAM2_OUT.awready,  -- out   std_logic;
            S_AXI_DRAM2_bresp    => S_AXI_DRAM2_OUT.bresp,    -- out   std_logic_vector(1 downto 0);
            S_AXI_DRAM2_bvalid   => S_AXI_DRAM2_OUT.bvalid,   -- out   std_logic;
            S_AXI_DRAM2_rdata    => S_AXI_DRAM2_OUT.rdata,    -- out   std_logic_vector(63 downto 0);
            S_AXI_DRAM2_rlast    => S_AXI_DRAM2_OUT.rlast,    -- out   std_logic;
            S_AXI_DRAM2_rresp    => S_AXI_DRAM2_OUT.rresp,    -- out   std_logic_vector(1 downto 0);
            S_AXI_DRAM2_rvalid   => S_AXI_DRAM2_OUT.rvalid,   -- out   std_logic;
            S_AXI_DRAM2_wready   => S_AXI_DRAM2_OUT.wready,   -- out   std_logic;
            S_AXI_DRAM3_araddr   => S_AXI_DRAM3_IN.araddr,    -- in    std_logic_vector(31 downto 0);
            S_AXI_DRAM3_arburst  => S_AXI_DRAM3_IN.arburst,   -- in    std_logic_vector(1 downto 0);
            S_AXI_DRAM3_arcache  => S_AXI_DRAM3_IN.arcache,   -- in    std_logic_vector(3 downto 0);
            S_AXI_DRAM3_arlen    => S_AXI_DRAM3_IN.arlen,     -- in    std_logic_vector(7 downto 0);
            S_AXI_DRAM3_arlock   => S_AXI_DRAM3_IN.arlock,    -- in    std_logic_vector(0 to 0);
            S_AXI_DRAM3_arprot   => S_AXI_DRAM3_IN.arprot,    -- in    std_logic_vector(2 downto 0);
            S_AXI_DRAM3_arqos    => S_AXI_DRAM3_IN.arqos,     -- in    std_logic_vector(3 downto 0);
            S_AXI_DRAM3_arregion => S_AXI_DRAM3_IN.arregion,  -- in    std_logic_vector(3 downto 0);
            S_AXI_DRAM3_arsize   => S_AXI_DRAM3_IN.arsize,    -- in    std_logic_vector(2 downto 0);
            S_AXI_DRAM3_arvalid  => S_AXI_DRAM3_IN.arvalid,   -- in    std_logic;
            S_AXI_DRAM3_awaddr   => S_AXI_DRAM3_IN.awaddr,    -- in    std_logic_vector(31 downto 0);
            S_AXI_DRAM3_awburst  => S_AXI_DRAM3_IN.awburst,   -- in    std_logic_vector(1 downto 0);
            S_AXI_DRAM3_awcache  => S_AXI_DRAM3_IN.awcache,   -- in    std_logic_vector(3 downto 0);
            S_AXI_DRAM3_awlen    => S_AXI_DRAM3_IN.awlen,     -- in    std_logic_vector(7 downto 0);
            S_AXI_DRAM3_awlock   => S_AXI_DRAM3_IN.awlock,    -- in    std_logic_vector(0 to 0);
            S_AXI_DRAM3_awprot   => S_AXI_DRAM3_IN.awprot,    -- in    std_logic_vector(2 downto 0);
            S_AXI_DRAM3_awqos    => S_AXI_DRAM3_IN.awqos,     -- in    std_logic_vector(3 downto 0);
            S_AXI_DRAM3_awregion => S_AXI_DRAM3_IN.awregion,  -- in    std_logic_vector(3 downto 0);
            S_AXI_DRAM3_awsize   => S_AXI_DRAM3_IN.awsize,    -- in    std_logic_vector(2 downto 0);
            S_AXI_DRAM3_awvalid  => S_AXI_DRAM3_IN.awvalid,   -- in    std_logic;
            S_AXI_DRAM3_bready   => S_AXI_DRAM3_IN.bready,    -- in    std_logic;
            S_AXI_DRAM3_rready   => S_AXI_DRAM3_IN.rready,    -- in    std_logic;
            S_AXI_DRAM3_wdata    => S_AXI_DRAM3_IN.wdata,     -- in    std_logic_vector(63 downto 0);
            S_AXI_DRAM3_wlast    => S_AXI_DRAM3_IN.wlast,     -- in    std_logic;
            S_AXI_DRAM3_wstrb    => S_AXI_DRAM3_IN.wstrb,     -- in    std_logic_vector(7 downto 0);
            S_AXI_DRAM3_wvalid   => S_AXI_DRAM3_IN.wvalid,    -- in    std_logic;
            S_AXI_DRAM3_arready  => S_AXI_DRAM3_OUT.arready,  -- out   std_logic;
            S_AXI_DRAM3_awready  => S_AXI_DRAM3_OUT.awready,  -- out   std_logic;
            S_AXI_DRAM3_bresp    => S_AXI_DRAM3_OUT.bresp,    -- out   std_logic_vector(1 downto 0);
            S_AXI_DRAM3_bvalid   => S_AXI_DRAM3_OUT.bvalid,   -- out   std_logic;
            S_AXI_DRAM3_rdata    => S_AXI_DRAM3_OUT.rdata,    -- out   std_logic_vector(63 downto 0);
            S_AXI_DRAM3_rlast    => S_AXI_DRAM3_OUT.rlast,    -- out   std_logic;
            S_AXI_DRAM3_rresp    => S_AXI_DRAM3_OUT.rresp,    -- out   std_logic_vector(1 downto 0);
            S_AXI_DRAM3_rvalid   => S_AXI_DRAM3_OUT.rvalid,   -- out   std_logic;
            S_AXI_DRAM3_wready   => S_AXI_DRAM3_OUT.wready    -- out   std_logic;
            );

end structural;